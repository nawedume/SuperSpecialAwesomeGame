
module collision_detector(
    input [4:0] current_x_pos,
    input [4:0] current_y_pos,
    input [2:0] move,
    input [1:0] map,
    input clk,
    output [4:0] new_x_pos,
    output [4:0] new_y_pos
);


        reg [19:0] i;
        always @(posedge clk) begin
            i <= i + 1;
        end
        always @(*) begin
            case(i) 
                20'd00: map1[0] = 20'b11111111011111111111;
                20'd01: map1[1] = 20'b10000001000100000001;
                20'd02: map1[2] = 20'b10000001000100000001;
                20'd03: map1[3] = 20'b10000001000100000001;
                20'd04: map1[4] = 20'b10000001000100000001;
                20'd05: map1[5] = 20'b10000000000100000001;
                20'd06: map1[6] = 20'b10000001111100011001;
                20'd07: map1[7] = 20'b10000000000000011001;
                20'd08: map1[8] = 20'b10000000000000011001;
                20'd09: map1[9] = 20'b11111111111111111001;
                20'd10: map1[10] = 20'b11111111111111111001;
                20'd11: map1[11] = 20'b11000000000000000001;
                20'd12: map1[12] = 20'b11000000000000000001;
                20'd13: map1[13] = 20'b11000000000000000001;
                20'd14: map1[14] = 20'b11111111111110111111;
            endcase
        end
        always @(*) begin
            case(i) 
                20'd00: map2[0] = 20'b11111111011111111111;
                20'd01: map2[1] = 20'b11111111010000000001;
                20'd02: map2[2] = 20'b11111111010000000001;
                20'd03: map2[3] = 20'b10000000010111111001;
                20'd04: map2[4] = 20'b10000000000000001001;
                20'd05: map2[5] = 20'b10111111111111111001;
                20'd06: map2[6] = 20'b10100000000100000001;
                20'd07: map2[7] = 20'b10100111100100000001;
                20'd08: map2[8] = 20'b10100100000100000001;
                20'd09: map2[9] = 20'b10100111111100000001;
                20'd10: map2[10] = 20'b10100000000000000001;
                20'd11: map2[11] = 20'b10111111111111111001;
                20'd12: map2[12] = 20'b10000000000010001001;
                20'd13: map2[13] = 20'b10000000000010001001;
                20'd14: map2[14] = 20'b11111111111110111111;
            endcase
        end
        always @(*) begin
            case(i) 
                20'd00: map3[0] = 20'b11111111011111111111;
                20'd01: map3[1] = 20'b11111111010000000001;
                20'd02: map3[2] = 20'b11111111010000000001;
                20'd03: map3[3] = 20'b10000000010111111001;
                20'd04: map3[4] = 20'b10000000000000001001;
                20'd05: map3[5] = 20'b10111111111111111001;
                20'd06: map3[6] = 20'b10100000000100000001;
                20'd07: map3[7] = 20'b10100111100100000001;
                20'd08: map3[8] = 20'b10100100000100000001;
                20'd09: map3[9] = 20'b10100111111100000001;
                20'd10: map3[10] = 20'b10100000000000000001;
                20'd11: map3[11] = 20'b10111111111111111001;
                20'd12: map3[12] = 20'b10000000000010001001;
                20'd13: map3[13] = 20'b10000000000010000001;
                20'd14: map3[14] = 20'b11111111111110111111;
            endcase
        end

    reg [0:19] current_map [0:14];
    reg [0:19] map1 [0:14];
    reg [0:19] map2 [0:14];
    reg [0:19] map3 [0:14];
    reg [0:19] map4 [0:14];

    // Draw maps here
    // MAP 1
    /*
    initial begin
        map1[0]     = 20'b11111111111111111111;
        map1[1]     = 20'b10000000000000000001;
        map1[2]     = 20'b10000000000000000001;
        map1[3]     = 20'b10000000000000000001;
        map1[4]     = 20'b10000000000000000001;
        map1[5]     = 20'b10000000000000000001;
        map1[6]     = 20'b10000000000000000001;
        map1[7]     = 20'b10000000000000000001;
        map1[8]     = 20'b10000000000000000001;
        map1[9]     = 20'b10000000000000000001;
        map1[10]    = 20'b10000000000000000001;
        map1[11]    = 20'b10000000000000000001;
        map1[12]    = 20'b10000000000000000001;
        map1[13]    = 20'b10000000000000000001;
        map1[14]    = 20'b11111111111111111111;
        map2[0]     = 20'b11111111111111111111;
        map2[1]     = 20'b10000000000000000001;
        map2[2]     = 20'b10000000000000000001;
        map2[3]     = 20'b10000000000000000001;
        map2[4]     = 20'b10000000000000000001;
        map2[5]     = 20'b10000000000000000001;
        map2[6]     = 20'b10000000000000000001;
        map2[7]     = 20'b10000000000000000001;
        map2[8]     = 20'b10000000000000000001;
        map2[9]     = 20'b10000000000000000001;
        map2[10]    = 20'b10000000000000000001;
        map2[11]    = 20'b10000000000000000001;
        map2[12]    = 20'b10000000000000000001;
        map2[13]    = 20'b10000000000000000001;
        map2[14]    = 20'b11111111111111111111;
        map3[0]     = 20'b11111111111111111111;
        map3[1]     = 20'b10000000000000000001;
        map3[2]     = 20'b10000000000000000001;
        map3[3]     = 20'b10000000000000000001;
        map3[4]     = 20'b10000000000000000001;
        map3[5]     = 20'b10000000000000000001;
        map3[6]     = 20'b10000000000000000001;
        map3[7]     = 20'b10000000000000000001;
        map3[8]     = 20'b10000000000000000001;
        map3[9]     = 20'b10000000000000000001;
        map3[10]    = 20'b10000000000000000001;
        map3[11]    = 20'b10000000000000000001;
        map3[12]    = 20'b10000000000000000001;
        map3[13]    = 20'b10000000000000000001;
        map3[14]    = 20'b11111111111111111111;
        map4[0]     = 20'b11111111111111111111;
        map4[1]     = 20'b10000000000000000001;
        map4[2]     = 20'b10000000000000000001;
        map4[3]     = 20'b10000000000000000001;
        map4[4]     = 20'b10000000000000000001;
        map4[5]     = 20'b10000000000000000001;
        map4[6]     = 20'b10000000000000000001;
        map4[7]     = 20'b10000000000000000001;
        map4[8]     = 20'b10000000000000000001;
        map4[9]     = 20'b10000000000000000001;
        map4[10]    = 20'b10000000000000000001;
        map4[11]    = 20'b10000000000000000001;
        map4[12]    = 20'b10000000000000000001;
        map4[13]    = 20'b10000000000000000001;
        map4[14]    = 20'b11111111111111111111;
    end
    */
    
    reg [4:0] temp_x;
    reg [4:0] temp_y;

    
    reg cc;

    
    always @ (*)
    begin

        if (move == 3'b100) begin   // RIGHT
                temp_x = current_x_pos + 1'b1;
                temp_y = current_y_pos;
            end
        
        else if (move == 3'b001) begin   // UP
                temp_x = current_x_pos;
                temp_y = current_y_pos - 1'b1;
            end
        
        else if (move == 3'b010) begin      // LEFT
                temp_x = current_x_pos - 1'b1;
                temp_y = current_y_pos;
            end
        
        else if (move == 3'b011) begin       // DOWN
                temp_x = current_x_pos;
                temp_y = current_y_pos + 1'b1;
            end
        
        else begin
            temp_x = current_x_pos;
            temp_y = current_y_pos;
        end

    end
    
    // Check if collision happened with new values
    always @ (move)
    begin
      case (map)
        2'b00: cc = map1[temp_x][temp_y];
        2'b01: cc = map2[temp_x][temp_y];
        2'b10: cc = map3[temp_x][temp_y];
        2'b11: cc = map4[temp_x][temp_y];
      endcase
    end


    // If collision happened retatin old value, if not go to new.
    assign new_x_pos = cc ? current_x_pos : temp_x;
    assign new_y_pos = cc ? current_y_pos : temp_y;
endmodule
